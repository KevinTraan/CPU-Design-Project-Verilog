//`include "gen_reg32_TB.svh"
//`include "mdr_TB.svh"
//`include "adder32_TB.svh"
//`include "sub32_TB.svh"
//`include "not32_TB.svh"
//`include "neg32_TB.svh"
//`include "ror32_TB.svh"
//`include "ShiftLeft_TB.svh"
`include "LAB_ROR_TB.svh"
//`include "LAB_SHR_TB.svh"
//`include "test_TB.svh"
//`include "DIV_TB.svh"