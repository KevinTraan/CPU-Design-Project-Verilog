`include "clock.svh"
`include "gen_reg32.svh"
`include "mux2to1.svh"
`include "mdr.svh"
`include "adder32.svh"
`include "adder16.svh"
`include "adder4.svh"
`include "sub32.svh"
`include "not32.svh"
`include "neg32.svh"
`include "ror32.svh"
`include "rol32.svh"
`include "Encoder_32_to_5.svh"
`include "Mux32to1.svh"
`include "bus.svh"
`include "ShiftLeft.svh"
`include "ShiftRight.svh"
`include "DIV.svh"
`include "ALU.svh"
`include "booth_mult.svh"