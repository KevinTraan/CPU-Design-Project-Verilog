`include "clock.svh"
`include "gen_reg32.svh"
`include "mux2to1.svh"
`include "mdr.svh"
`include "Encoder_32_to_5.svh"
`include "Mux32to1.svh"
`include "bus.svh"
`include "ALU.svh"
`include "reg0.svh"
`include "con_FF.svh"
`include "MAR_RAM.svh"
`include "select_logic.svh"
`include "pc_reg.svh"
`include "ra.svh"
`include "In_Port.svh"
